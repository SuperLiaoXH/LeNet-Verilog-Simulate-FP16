// ----------------------------------------------------------------------------------
// -- Function : This module is the design of LeNet-5
// -- Designer : LXH
// ----------------------------------------------------------------------------------
module LeNet
(

);


endmodule